//module
//endmodule
