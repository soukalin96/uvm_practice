//module 

//endmodule
