//module
//edit 1
//endmodule
